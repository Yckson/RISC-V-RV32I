
module Plus4 (
    input wire [63:0] PC,
    output wire [63:0] Plus4
);
    
endmodule

assign Plus4 = PC + 4;